`timescale 1ns / 1ns

module scoreboard(

    );
endmodule
