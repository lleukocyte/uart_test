`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.08.2025 19:56:07
// Design Name: 
// Module Name: environment
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

class env extends uvm_env;
    `uvm_component_utils(env);
    
   sequencer sequencer_h;
   driver driver_h;
   monitor monitor_h;
   scoreboard scoreboard_h;
   monitor monitor_h;
   
   function new (string name, uvm_component parent);
      super.new(name,parent);
   endfunction : new

   function void build_phase(uvm_phase phase);
      sequencer_h = new("sequencer_h",this);
      driver_h = driver::type_id::create("driver_h",this);
      monitor_h = monitor::type_id::create("monitor_h",this);
      coverage_h    = coverage::type_id::create ("coverage_h",this);
      scoreboard_h  = scoreboard::type_id::create("scoreboard",this);
   endfunction : build_phase

   function void connect_phase(uvm_phase phase);

      driver_h.seq_item_port.connect(sequencer_h.seq_item_export);

      monitor_h.ap.connect(coverage_h.analysis_export);
      monitor_h.ap.connect(scoreboard_h.data_f.analysis_export);
   endfunction : connect_phase
endclass