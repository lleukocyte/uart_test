`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/26/2025 02:23:39 PM
// Design Name: 
// Module Name: test_pkg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


package test_pkg;
    `include "sequence_item.sv"
    `include "sequence.sv"
    `include "sequencer.sv"
    `include "scoreboard.sv"
    `include "monitor.sv"
    `include "driver.sv"
    `include "agent.sv"
    `include "environment.sv"
    `include "base_test.sv"
endpackage